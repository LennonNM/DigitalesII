module NAND ();

  





endmodule
